library verilog;
use verilog.vl_types.all;
entity Group_16_vlg_vec_tst is
end Group_16_vlg_vec_tst;
