-- ELECTENG 209 UART_ Receiver
-- Last Edit: 2016/08/12

-------------------------------------------------------
-----------            S Counter            -----------
-------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity s_counter is
	port (
		clk, reset_S	:	in	std_logic;
		enable_S			:	in std_logic;
		s_cnt 			:	buffer std_logic_vector(3 downto 0));
end entity;

architecture beh of s_counter is
begin
	process (clk, reset_S)
		begin
			if rising_edge(clk) then
				if reset_S = '1' then
					s_cnt <= B"0000";
				elsif (reset_S	= '0' AND enable_S = '1') then
					s_cnt <= s_cnt + 1;
				end if;
			end if;
	end process;
end beh;

-------------------------------------------------------
-----------            N Counter            -----------
-------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity n_counter is
	port (
		clk, reset_N	:	in	std_logic;
		enable_N			:	in std_logic;
		n_cnt 			:	buffer std_logic_vector(3 downto 0));
end entity;

architecture beh of n_counter is
begin
	process (clk, reset_N)
		begin
			if rising_edge(clk) then
				if reset_N = '1' then
					n_cnt <= B"0000";
				elsif (reset_N	= '0' AND enable_N = '1') then
					n_cnt <= n_cnt + 1;
				end if;
			end if;
	end process;
end beh;

-------------------------------------------------------
-----------         S Comparator 7          -----------
-------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity s_comp_7 is
	port (
		s_cnt 			:	in std_logic_vector(3 downto 0);
		cmp7_s			:	out std_logic);		
end entity;

architecture beh of s_comp_7 is
begin
	process (s_cnt)
		begin
			if s_cnt = B"0111" then
				cmp7_s <= '1';
			else
				cmp7_s <= '0';
			end if;
	end process;
end beh;


-------------------------------------------------------
-----------        S Comparator 15          -----------
-------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity s_comp_15 is
	port (
		s_cnt 			:	in std_logic_vector(3 downto 0);
		cmp15_s			:	out std_logic);		
end entity;

architecture beh of s_comp_15 is
begin
	process (s_cnt)
		begin
			if s_cnt = B"1111" then
				cmp15_s <= '1';
			else
				cmp15_s <= '0';
			end if;
	end process;
end beh;

-------------------------------------------------------
-----------         N Comparator 7          -----------
-------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity n_comp_7 is
	port (
		n_cnt 			:	in std_logic_vector(3 downto 0);
		cmp7_n			:	out std_logic);		
end entity;

architecture beh of n_comp_7 is
begin
	process (n_cnt)
		begin
			if n_cnt = B"0111" then
				cmp7_n <= '1';
			else
				cmp7_n <= '0';
			end if;
	end process;
end beh;

-------------------------------------------------------
-----------         Shift Register          -----------
-------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity shift_reg is
	port (
		clk, enable_shift, rx:	in std_logic;
		buf	: buffer std_logic_vector(7 DOWNTO 0));	
end entity;

architecture beh of shift_reg is 
begin
	process (clk)
		begin
			if rising_edge(clk) then
				if enable_shift = '1' then
					buf(7 DOWNTO 0) <= rx & buf(7 DOWNTO 1);
				end if;
			end if;
	end process;
end beh;

-------------------------------------------------------
-----------             BCD2SSD             -----------
-------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity BCD2SSD is
port(
	clk : in std_logic;
	bcd : in std_logic_vector(7 downto 0);
	segment7 : out std_logic_vector(6 downto 0);
	decptn	:	out std_logic;
	digit : out std_logic_vector(3 downto 0));
end BCD2SSD;

architecture beh of BCD2SSD is
	signal SEG : std_logic_vector(1 downto 0);
	signal DIS : std_logic_vector(3 downto 0);
begin
	process (clk,bcd)
		begin
			SEG(1 downto 0) <= bcd(6 downto 5);
			DIS(3 downto 0) <= bcd(3 downto 0);
			if rising_edge(clk) then
				decptn <= bcd(4);
				case SEG is
					when "00"=> digit <="0001";
					when "01"=> digit <="0010";
					when "10"=> digit <="0100";
					when "11"=> digit <="1000";
					when others=> digit <="0000";
				end case;
				case DIS is
					when "0000"=> segment7 <="0111111";
					when "0001"=> segment7 <="0000110";
					when "0010"=> segment7 <="1011011";
					when "0011"=> segment7 <="1001111";
					when "0100"=> segment7 <="1100110";
					when "0101"=> segment7 <="1101101";
					when "0110"=> segment7 <="1111101";
					when "0111"=> segment7 <="0000111";
					when "1000"=> segment7 <="1111111";
					when "1001"=> segment7 <="1101111";
					when "1010"=> segment7 <="1110111";
					when "1011"=> segment7 <="1111100";
					when "1100"=> segment7 <="0111001";
					when "1101"=> segment7 <="1011110";
					when "1110"=> segment7 <="1111011";
					when "1111"=> segment7 <="1110001";
					when others=> segment7 <="0000000";
				end case;
			end if;
	end process;
end beh;

-------------------------------------------------------
-----------            Register             -----------
-------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity parallel_register is
port(
	parallel_in : in std_logic_vector(7 downto 0);
	load, clk : in std_logic;
	parallel_out: out std_logic_vector(7 downto 0)
); end parallel_register;

architecture beh of parallel_register is 

begin
	process (clk)
	begin
		if rising_edge(clk) then
			if load = '1' then
				parallel_out <= parallel_in;
			end if;	
		end if;
	end process;
end beh;	

------------------------------------------------------
------------------- Counter 2 ------------------------
------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Counter2_VHDL is
   port(clk: in std_logic;
		  bcd_out: out std_logic_vector(7 downto 0));
end Counter2_VHDL;

architecture beh of Counter2_VHDL is
   signal temp: std_logic_vector(7 downto 0);
begin
	process(clk)
   begin
      if rising_edge(clk) then
			case temp is
				when x"00"=> bcd_out <=x"6E";
				when x"01"=> bcd_out <=x"4A";
				when x"02"=> bcd_out <=x"3A";
				when others=> bcd_out <=x"00";
			end case;
			if temp=x"02" then
				temp<=x"00";
			else
				temp <= temp + 1;
			end if;
      end if;
   end process;
end beh;

-------------------------------------------------------
-----------               MUX               -----------
-------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity mux is
	port (
		idle			:	in	std_logic;
		ina,inb		:	in std_logic_vector(7 downto 0);
		bcd_out		: out std_logic_vector(7 downto 0));
end entity;


architecture beh of mux is
begin
	with idle select bcd_out <= ina when '0', inb when '1';
end architecture;

-------------------------------------------------------
-----------               FSM               -----------
-------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity fsm is
	port (
		clk			:	in	std_logic;
		rx				:	in std_logic;
		reset_N, reset_S, enable_N, enable_S, enable_shift, load, sid : out std_logic;
		cmp15_s, cmp7_s, cmp7_n : in std_logic);
end entity;

--Define architecture here 

architecture beh of fsm is

	type my_states is (idle, start, data, stop,finish);
	signal CS, NS : my_states:= idle;

begin

	----------------------------
	--VHDL code for FSM
	----------------------------

	--state registers
	Synchronous_process: process (clk)
		begin
			if rising_edge(clk) then
				CS <= NS;
			end if;
	end process;
			
	------------------------------------

	NextState_logic: process (CS, rx, cmp15_s, cmp7_n, cmp7_s)
		begin
			case CS is
				when idle =>
					if rx = '0' then
						NS <= start;
					else
						NS <= idle;
					end if;
				when start =>
					if (cmp7_s = '1' AND rx = '0') then
						NS <= data;
					elsif cmp15_s = '1' then
						NS <= idle;
					else
						NS <= start;
					end if;
				when data =>
					if (cmp15_s = '1' AND cmp7_n = '1') then
						NS <= stop;
					else
						NS <= data;
					end if;
				when stop =>
					if cmp15_s = '0' then
						NS <= stop;
					else
						NS <= finish;
					end if;
				when finish =>
					if cmp7_s = '1' then
						NS <= idle;
					else
						NS <= finish;
					end if;
			end case;
	end process;

	-----------------------------------------

	Output_logic: process (CS, rx, cmp15_s, cmp7_n, cmp7_s)
		begin
		enable_shift <= '0';
		reset_S <= '0';
		reset_N <= '0';
		enable_N <= '0';
		enable_S <= '0';
		load <= '0';
			case CS is
				when idle =>
					if rx = '0' then
						reset_S <= '1';
					else
						reset_S <= '0';
					end if;
					sid <= '1';
				when start =>
					if cmp7_s = '1' then
						reset_S <= '1';
						reset_N <= '1';
					elsif (cmp15_s = '1') then
						reset_S <= '1';
					else
						enable_S <= '1';
					end if;
					sid <= '0';
				when data =>
					if (cmp7_n = '1' AND cmp15_s = '1') then
						reset_S <= '1';
						enable_shift <= '1';
					elsif (cmp7_n = '0' AND cmp15_s = '1') then
						enable_shift <= '1';
						reset_S <= '1';
						enable_N <= '1';
					else
						enable_S <= '1';
					end if;
					sid <= '0';
				when stop =>
					if cmp15_s = '0' then
						enable_S <= '1';
					else
						enable_S <= '0';
					end if;
					sid <= '0';
				when finish =>
					if cmp7_s = '1' then
						load <= '1';
					else
						enable_S <= '1';
					end if;
					sid <= '0';
			end case;
	end process;
end beh;